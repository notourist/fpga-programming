module ascon();
endmodule
