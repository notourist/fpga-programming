module gpio();
endmodule
